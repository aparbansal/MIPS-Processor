module processor();

endmodule
